-------------------------------------------------------------------------
--Christopher hausner & Caden Otis
-- Iowa State University
-------------------------------------------------------------------------


-- Fiveto32Decoder.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of a Fiveto32Decoder
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity Fiveto32Decoder is

  port(i_EN          : in std_logic;
       i_D          : in std_logic_vector(4 downto 0);
       o_O          : out std_logic_vector(31 downto 0));

end Fiveto32Decoder;

architecture dataflow of Fiveto32Decoder is
begin
		  o_O <=    "00000000000000000000000000000001" when (i_D = "00000" and i_EN = '1') else
					"00000000000000000000000000000010" when (i_D = "00001" and i_EN = '1') else
					"00000000000000000000000000000100" when (i_D = "00010" and i_EN = '1') else
					"00000000000000000000000000001000" when (i_D = "00011" and i_EN = '1') else
					"00000000000000000000000000010000" when (i_D = "00100" and i_EN = '1') else
					"00000000000000000000000000100000" when (i_D = "00101" and i_EN = '1') else
					"00000000000000000000000001000000" when (i_D = "00110" and i_EN = '1') else
					"00000000000000000000000010000000" when (i_D = "00111" and i_EN = '1') else
					"00000000000000000000000100000000" when (i_D = "01000" and i_EN = '1') else
					"00000000000000000000001000000000" when (i_D = "01001" and i_EN = '1') else
					"00000000000000000000010000000000" when (i_D = "01010" and i_EN = '1') else
					"00000000000000000000100000000000" when (i_D = "01011" and i_EN = '1') else
					"00000000000000000001000000000000" when (i_D = "01100" and i_EN = '1') else
					"00000000000000000010000000000000" when (i_D = "01101" and i_EN = '1') else
					"00000000000000000100000000000000" when (i_D = "01110" and i_EN = '1') else
					"00000000000000001000000000000000" when (i_D = "01111" and i_EN = '1') else
					"00000000000000010000000000000000" when (i_D = "10000" and i_EN = '1') else
					"00000000000000100000000000000000" when (i_D = "10001" and i_EN = '1') else
					"00000000000001000000000000000000" when (i_D = "10010" and i_EN = '1') else
					"00000000000010000000000000000000" when (i_D = "10011" and i_EN = '1') else
					"00000000000100000000000000000000" when (i_D = "10100" and i_EN = '1') else
					"00000000001000000000000000000000" when (i_D = "10101" and i_EN = '1') else
					"00000000010000000000000000000000" when (i_D = "10110" and i_EN = '1') else
					"00000000100000000000000000000000" when (i_D = "10111" and i_EN = '1') else
					"00000001000000000000000000000000" when (i_D = "11000" and i_EN = '1') else
					"00000010000000000000000000000000" when (i_D = "11001" and i_EN = '1') else
					"00000100000000000000000000000000" when (i_D = "11010" and i_EN = '1') else
					"00001000000000000000000000000000" when (i_D = "11011" and i_EN = '1') else
					"00010000000000000000000000000000" when (i_D = "11100" and i_EN = '1') else
					"00100000000000000000000000000000" when (i_D = "11101" and i_EN = '1') else
					"01000000000000000000000000000000" when (i_D = "11110" and i_EN = '1') else
					"10000000000000000000000000000000" when (i_D = "11111" and i_EN = '1') else
					(others => '0');
end dataflow;
